//////////////////////////////////////////////////////////////////////////////////
// Engineer: Yurin VV
// Create Date: 07.2022
// Module Name: parameters
// Project Name: Some DAC
// Tool Versions: Vivado 2018.2
// Description: Offsets in a register group
//////////////////////////////////////////////////////////////////////////////////	parameter LINEA_OFFSET   = 0;
parameter LINET_OFFSET   = 9;
parameter LINENMB_OFFSET = 18;
parameter REPEATCYCLE    = 19;
parameter INC_OFFSET     = 20;
parameter END_OFFSET     = 28;
parameter LINET_F_OFFSET = 29;
parameter LINET_F_END    = 38;